module i2s_rx (
);

endmodule
