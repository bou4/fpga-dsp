module i2s_rx (
);

    // TODO

endmodule
